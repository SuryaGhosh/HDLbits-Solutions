module top_module ( 
    input [15:0] a, b,
    input cin,
    output cout,
    output [15:0] sum );
    wire [0:0] cout_1, cout_2, cout_3; 
    
    bcd_fadd fadd1(.a(a[3:0]), .b(b[3:0]), .cin(cin), .cout(cout_1), .sum(sum[3:0]));
    bcd_fadd fadd2(.a(a[7:4]), .b(b[7:4]), .cin(cout_1), .cout(cout_2), .sum(sum[7:4]));
    bcd_fadd fadd3(.a(a[11:8]), .b(b[11:8]), .cin(cout_2), .cout(cout_3), .sum(sum[11:8]));    
    bcd_fadd fadd4(.a(a[15:12]), .b(b[15:12]), .cin(cout_3), .cout(cout), .sum(sum[15:12]));
endmodule


