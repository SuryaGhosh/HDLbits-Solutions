module top_module (
    input clk,
    input reset,
    output OneHertz,
    output [2:0] c_enable
); 
    
    // 1 cycle/second = 1 hz
    // divide the input signal by 10, 3 times 
    // we have 3 chained counters, each counter counts to 10
    wire [3:0] Q0, Q1, Q2;
    
    assign OneHertz = (Q2 == 4'b1001 & Q1 == 4'b1001 & Q0 == 4'b1001);
    assign c_enable[0] = 1'b1;
    assign c_enable[1] = (Q0 == 4'b1001);
    assign c_enable[2] = (Q0 == 4'b1001 & Q1 == 4'b1001);
    
    bcdcount counter0 (.clk(clk), .reset(reset), .enable(c_enable[0]), .Q(Q0));
    bcdcount counter1 (.clk(clk), .reset(reset), .enable(c_enable[1]), .Q(Q1));
    bcdcount counter2 (.clk(clk), .reset(reset), .enable(c_enable[2]), .Q(Q2));

endmodule

